library ieee;
use ieee.std_logic_1164.all;

entity multi_barrel_testing is
    